//--------------------------------------------------
// Created by : Teodor Dimitrov
// Design     : async_fifo
// Module name: async_fifo_sequencer.sv
//
// Description: UVM sequencer for the async FIFO module.
//              Extends uvm_sequencer class
//




